{
"project_title": "INTELLIGENT BEDÖMNING AV RISKNIVÅER FÖR ALLVARA ARRHYTHMIAS",
"h1_credits": "Uppskattning av risknivån för arytmi",
"h2_credits": "Projektkrediter",
"h1_login": "Arytmi risk nivå",
"h2_login": "Logga in",
"h3_login": "Medarbetare",
"login": "Logga in",
"university": "Jaens Universitet",
"quiron": "Hospital Universitario QuirónSalud de Madrid",
"sas": "Complejo Hospitalario de Jaén y Linares",
"avs": "Hospital General Universitario de Elda",
"h1_menu": "Arytmi risk nivå  ",
"ecg": "ECG",
"ecg_done": "ECG Genomförda",
"patients": "Patienter",
"logout": "Logga ut",
"return": "Gå tillbaka",
"h1_logout": "Logga ut",
"h2_logout": "Är du säker på att du vill logga ut?",
"accept": "Acceptera",
"deny": "Avbryt",
"h1_record": "Historik ECG",
"h2_record": "Historik ECG",
"search": "Söka efter",
"dni": "Identifierare",
"date": "Datum",
"risklevel": "Risk nivå",
"riskcontext": "Klinik information",
"actions": "Vidtagna åtgärder",
"years": "År",
"male": "Man",
"female": "Kvinna",
"action1": "Öka frekvensen",
"action2": "Minska frekvensen",
"action3": "Granska behandlingen",
"action4": "Mätning 4",
"action5": "Mätning 5",
"riskfactor1": "Mer än 67",
"riskfactor2": "Kvinna",
"riskfactor3": "Diuretikum",
"riskfactor4": "Serum",
"riskfactor5": "Akut hjärtinfarkt",
"riskfactor6": "Sepsis",
"riskfactor7": "Ett läkemedel förlänger QT",
"riskfactor8": "Två eller fler läkemedel förlänger QT",
"riskfactor9": "Hjärt",
"tag_yes": "Ja ",
"tag_no": "Nej",
"h1_patients": "Patienter",
"h2_patients": "Ny/Uppdatera patienter",
"save": "Spara",
"name": "Namn",
"surname": "Efternamn",
"birthday": "Födelsedag",
"sex": "Kön",
"iam_label": "Akut hjärtinfarkt",
"cardiac_label": "Hjärtsvikt",
"remarks": "Anmärkningar",
"h1_ecg": "ECG",
"h2_ecg": "Arytmi risk nivå bedömning",
"estimate": "Beräkna",
"factors": "Faktorer",
"factor1": "Diuretikum ASA (furosemid, torasemide, bumetanid)",
"factor2": "Serum med kalium (K+) <=3,5 mEq/L",
"factor3": "Sepsis",
"factor4": "Ett läkemedel förlänger QT",
"factor5": "Två eller fler läkemedel förlänger QT",
"factors_legend": "Låg: 0 till 1.58 | Mellan: 1.59 till 2.38 | Hög: 2.39 till 5 ",
"risk": "Risk",
"risk_label":  "Odefinierad klinik information",
"risk_string": "Klinik information ",
"risk_undefined": "Odefinierad",
"risk_low": "Låg",
"risk_average": "Mellan",
"risk_high": "Hög",
"page": "Sida",
"next": "Nästa",
"prev": "Tidigare",
"prep": " Av ",
"iderror": "Där är ingen information om denna patienten!",
"notexist": "Patienten existerar inte!",
"computing": "Beräknad",
"qtcerror": "Kan inte beräkna QTc!",
"link2menu": "Meny",
"fileerror": "Ingen fil är vald!",
"exterror": "Fel förlängning",
"edit": "Redigera",
"basal_tx": "Basal",
"upfile1": "Lägg till ECG-bild",
"deletefile1": "Ta bort ECG-bild",
"clipped": "Ursprunglig klippning",
"qtc_man": "Ange värde, om tillgängligt",
"historial": "Patientens historia",
"actualiza": "Uppdatera observationer",
"number": "Siffra",
"actualizaecg": "Uppdatera och gå tillbaka till historiken"
}